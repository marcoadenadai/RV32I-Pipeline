LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;

ENTITY MUX_ALU_1 IS
   PORT (
		BRANCH_DO_IT: IN STD_LOGIC;
		PC_IN_MUX		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		REG_OUT_1	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		MUX_OUT_ALU_1	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
END ENTITY;

ARCHITECTURE MUX_ALU_1_Arch OF MUX_ALU_1 IS
	
	BEGIN
		WITH BRANCH_DO_IT SELECT 
		   MUX_OUT_ALU_1 <= PC_IN_MUX WHEN '1',
								  REG_OUT_1 WHEN '0',
								  REG_OUT_1 WHEN OTHERS;
								  

		
END ARCHITECTURE;