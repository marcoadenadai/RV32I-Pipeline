LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE REGPIPE_ID_EX_PACKAGE IS
   COMPONENT REGPIPE_ID_EX 
   PORT (
      clock    				: IN STD_LOGIC := '0';
		Reset						: IN STD_LOGIC := '0';
		PCIn						: IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
      PCOut        			: OUT STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
		REG_1_IN       		: IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
      REG_1_OUT		      : OUT STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
		REG_2_IN       		: IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
      REG_2_OUT			   : OUT STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
		InstructionIn			: IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
      InstructionOut       : OUT STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
		
		ctl_RegWrite_IN		: IN STD_LOGIC := '0';
		ctl_RegWrite_OUT		: OUT STD_LOGIC := '0';
		
		ctl_MemToReg_IN		: IN STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
		ctl_MemToReg_OUT		: OUT STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
		
		ctl_MemWrite_IN		: IN STD_LOGIC := '0';
		ctl_MemWrite_OUT		: OUT STD_LOGIC := '0';
		
		ctl_MemRead_IN			: IN STD_LOGIC := '0';
		ctl_MemRead_OUT		: OUT STD_LOGIC := '0';
		
		ctl_BranchDoIt_IN		: IN STD_LOGIC := '0';
		ctl_BranchDoIt_OUT	: OUT STD_LOGIC := '0';
		
		ctl_BranchOP_IN		: IN STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";
		ctl_BranchOP_OUT		: OUT STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";
		
		ctl_ALUSrc_IN			: IN STD_LOGIC := '0';
		ctl_ALUSrc_OUT			: OUT STD_LOGIC := '0';
		
		ctl_ALUOp_IN			: IN STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
		ctl_ALUOp_OUT			: OUT STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
		
		ctl_ImmType_IN			: IN STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";
		ctl_ImmType_OUT		: OUT STD_LOGIC_VECTOR(2 DOWNTO 0) := "000"
	);
   END COMPONENT;
END REGPIPE_ID_EX_PACKAGE;