LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE MUX_ALU_1_PACKAGE IS
   COMPONENT MUX_ALU_1
      PORT (
		BRANCH_DO_IT: IN STD_LOGIC;
		PC_IN_MUX		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		REG_OUT_1	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		MUX_OUT_ALU_1	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
   END COMPONENT;
END MUX_ALU_1_PACKAGE;