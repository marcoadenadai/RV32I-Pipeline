LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;

ENTITY PC_MUX IS
   PORT (
		BRANCH_CONTROL: IN STD_LOGIC;
		MUX_IN		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		BRANCH_IN	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		MUX_OUT	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
END ENTITY;

ARCHITECTURE PC_MUX_Arch OF PC_MUX IS
	
	BEGIN

      PROCESS (BRANCH_CONTROL)
      BEGIN
		
         IF BRANCH_CONTROL = '1' THEN
				MUX_OUT <= BRANCH_IN;
			ELSE
				MUX_OUT <= MUX_IN;		
         END IF;
			
      END PROCESS;
		
END ARCHITECTURE;