LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;

ENTITY REGPIPE_ID_EX IS
   PORT (
      clock    				: IN STD_LOGIC := '0';
		Reset						: IN STD_LOGIC := '0';
		PCIn						: IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
      PCOut        			: OUT STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
		REG_1_IN       		: IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
      REG_1_OUT		      : OUT STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
		REG_2_IN       		: IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
      REG_2_OUT			   : OUT STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
		InstructionIn			: IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
      InstructionOut       : OUT STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000"
		);
END ENTITY;

ARCHITECTURE REGPIPE_ID_EX_Arch OF REGPIPE_ID_EX IS
	BEGIN
      PROCESS (clock)
      BEGIN
		
         IF rising_edge(clock) THEN
				
				IF Reset = '1' THEN
					PCOut <= "00000000000000000000000000000000";
					InstructionOut <= "00000000000000000000000000000000";
					REG_1_OUT <= "00000000000000000000000000000000";
					REG_2_OUT <= "00000000000000000000000000000000";
				ELSE
					PCOut <= PcIn;
					REG_1_OUT <= REG_1_IN;
					REG_2_OUT <= REG_2_IN;
					InstructionOut <= InstructionIn;
				END IF;
				
         END IF;
			
      END PROCESS;
END ARCHITECTURE;