LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
use ieee.numeric_std.all;

ENTITY BRANCH_COMPARE IS
   PORT (
      clock    				: IN STD_LOGIC := '0';
		Reset						: IN STD_LOGIC := '0';
		BRANCH_OP				: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		REG_1_IN       		: IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
		REG_2_IN       		: IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
      DECISION       : OUT STD_LOGIC := '0'
		);
END ENTITY;

ARCHITECTURE BRANCH_COMPARE_Arch OF BRANCH_COMPARE IS
	
	SIGNAL SUB_S  : SIGNED(31 DOWNTO 0);
	SIGNAL SUB_U  : UNSIGNED(31 DOWNTO 0);
	
	--SIGNAL OP1_UNS  : unsigned(31 DOWNTO 0);
	--SIGNAL OP2_UNS  : unsigned(31 DOWNTO 0);
	
	
	
	BEGIN
      PROCESS (BRANCH_OP, REG_1_IN, REG_2_IN)
      BEGIN
			CASE BRANCH_OP IS
				WHEN "000" => 
				-- BEQ
						SUB_S <= SIGNED(REG_1_IN) - SIGNED(REG_2_IN);
						IF SUB_S = "000000000000000000000000000000" THEN 
							DECISION <= '1';
						ELSE 
							DECISION <= '0';
						END IF;
						 
				
				WHEN "001" =>
				-- BNE
						SUB_S <= SIGNED(REG_1_IN) - SIGNED(REG_2_IN);
						IF SUB_S = "000000000000000000000000000000" THEN 
							DECISION <= '0';
						ELSE 
							DECISION <= '1';
						END IF;
				
				
				WHEN "100" =>
				-- BLT
						SUB_S <= SIGNED(REG_1_IN) - SIGNED(REG_2_IN);
						IF SUB_S < "000000000000000000000000000000" THEN 
							DECISION <= '1';
						ELSE 
							DECISION <= '0';
						END IF;
				
				WHEN "101" =>
				-- BGE
						SUB_S <= SIGNED(REG_1_IN) - SIGNED(REG_2_IN);
						IF SUB_S > "000000000000000000000000000000" OR SUB_S = "000000000000000000000000000000" THEN 
							DECISION <= '1';
						ELSE 
							DECISION <= '0';
						END IF;
				
				WHEN "110" =>
				-- BLTU
						--OP1_UNS <= unsigned(REG_1_IN);
						--OP2_UNS <= unsigned(REG_2_IN);
						SUB_U <= UNSIGNED(REG_1_IN) - UNSIGNED(REG_2_IN);
						IF SUB_U < "000000000000000000000000000000" THEN 
							DECISION <= '1';
						ELSE 
							DECISION <= '0';
						END IF;
						
				
				WHEN "111" =>
				-- BGEU
						SUB_U <= UNSIGNED(REG_1_IN) - UNSIGNED(REG_2_IN);
						IF SUB_U > "000000000000000000000000000000" OR SUB_S = "000000000000000000000000000000" THEN 
							DECISION <= '1';
						ELSE 
							DECISION <= '0';
						END IF;
				
				WHEN OTHERS => NULL;
			
			END CASE;
      END PROCESS;
END ARCHITECTURE;

