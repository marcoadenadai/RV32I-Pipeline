LIBRARY ieee;
USE ieee.std_logic_1164.all;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY ADDER IS
    PORT (
        A	: IN STD_LOGIC_VECTOR (31 DOWNTO 0) := "00000000000000000000000000000000";
        S 	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0) := "00000000000000000000000000000000"
    );
END ENTITY;

ARCHITECTURE ADDER_arch OF ADDER IS
BEGIN
	S <= A + "00000000000000000000000000000001";
END ARCHITECTURE; 