LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE IMM_HANDLER_PACKAGE IS
   COMPONENT IMM_HANDLER
      PORT (
			IMM_TYPE				: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			INSTRUCTION       : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
			RD       		   : OUT STD_LOGIC_VECTOR(4 DOWNTO 0);
			IMM_OUT           : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
   END COMPONENT;
END IMM_HANDLER_PACKAGE;