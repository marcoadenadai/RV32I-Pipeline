LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE MUX_PC_PACKAGE IS
   COMPONENT PC_MUX 
   PORT (
      BRANCH_CONTROL: IN STD_LOGIC;
		MUX_IN		: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		BRANCH_IN	: IN STD_LOGIC_VECTOR(31 DOWNTO 0);
		MUX_OUT	: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);
   END COMPONENT;
END MUX_PC_PACKAGE;