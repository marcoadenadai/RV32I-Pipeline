LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;
USE ieee.std_logic_signed.all;

PACKAGE RAM_PACKAGE IS
   COMPONENT RAM
      PORT (
			CLOCK			: IN STD_LOGIC;
		  RESET			: IN STD_LOGIC;
		  MEM_WRITE    : IN STD_LOGIC;
		  MEM_READ		: IN STD_LOGIC;
        ADDR			: IN UNSIGNED(31 DOWNTO 0);
		  WRITE_DATA   : IN STD_LOGIC_VECTOR(31 DOWNTO 0);	
        MEM_OUT		: OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
   END COMPONENT;
END RAM_PACKAGE;