LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY work;
USE work.PC_PACKAGE.all;

USE work.ROM_PACKAGE.all;

USE work.REGPIPE_IF_DF_PACKAGE.all;

ENTITY PROCESSADOR IS
	PORT(
		CLK : IN STD_LOGIC;
		RESET: IN STD_LOGIC
		
		--Saida_PC : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		--Saida_ROM : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		--Saida_TEST : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);

END ENTITY;

ARCHITECTURE PROCESSADOR_ARCH OF PROCESSADOR IS
	--variable PC_IN: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL PC_OUT: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL PC_NEXT: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ROM_INSTRUCTION: STD_LOGIC_VECTOR(31 DOWNTO 0);


--	SIGNAL ROM_INSTRUCTION: STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
--	--SIGNAL TEST_RETURN: STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
--	SIGNAL REGPIPE_IF_DF_SAIDA_PC:  STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000"; --Serão as entrada do estágio de DF
--	SIGNAL REGPIPE_IF_DF_SAIDA_INSTRUCTION:  STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";--Serão as entrada do estágio de DF
--	
	SIGNAL myCLK: STD_LOGIC;
	SIGNAL myRESET: STD_LOGIC;
	
	
 BEGIN
	
	myCLK <= CLK;
	myRESET <= RESET;
 
	PC_C0: PC PORT MAP(myCLK, myRESET, PC_NEXT, PC_OUT, PC_NEXT);
	ROM_C1: ROM PORT MAP(myCLK, myRESET, PC_OUT, ROM_INSTRUCTION);
	

--	ROM_C1: ROM PORT MAP(PC_VALUE, ROM_INSTRUCTION, myCLK, myRESET);
--	
--	REGPIPE_IF_DF_C3: REGPIPE_IF_DF PORT MAP(myCLK, myRESET, PC_VALUE, REGPIPE_IF_DF_SAIDA_PC, ROM_INSTRUCTION, REGPIPE_IF_DF_SAIDA_INSTRUCTION);
--	
--	Saida_TEST <= REGPIPE_IF_DF_SAIDA_INSTRUCTION;
--	Saida_PC <= PC_VALUE;
--	Saida_ROM <= ROM_INSTRUCTION;
	
END ARCHITECTURE;