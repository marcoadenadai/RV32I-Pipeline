LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY ROM IS
    PORT (
		clock    : IN STD_LOGIC := '0';
		Reset 	: IN STD_LOGIC := '0';
      ADDR 		: IN STD_LOGIC_VECTOR (31 DOWNTO 0); -- ENDERECO DA MEMORIA DE INSTRUCAO 
      S 			: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
    );
END ENTITY;

ARCHITECTURE ROM_arch OF ROM IS

	signal fio_addr : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
	signal fio_result : std_logic_vector(31 downto 0);
	
	
BEGIN	
	fio_addr <= ADDR;
	S <= fio_result;
		
--		PROCESS (clock, Reset, fio_result)
--			variable var : std_logic_vector(31 downto 0);
--      BEGIN
--         IF rising_edge(clock) and Reset = '1' THEN
--					-- no momento de reset eu jogo a primeira instrucao que comeca a ROM
--					var := "00000000000000000000010110010011";
--					fio_result <= var;
--         END IF;
--			
--      END PROCESS;
	
		PROCESS (ADDR, clock) BEGIN --fio_addr
				CASE fio_addr IS
					WHEN "00000000000000000000000000000000" => fio_result <= "00000000000000000000010110010011";
					WHEN "00000000000000000000000000000001" => fio_result <= "00000000101000000000010100010011";
					WHEN "00000000000000000000000000000010" => fio_result <= "00000001000000000000000011101111";
					WHEN "00000000000000000000000000000011" => fio_result <= "00000001111000000000010100010011";
					WHEN "00000000000000000000000000000100" => fio_result <= "00000001111100000000010100010011";
					WHEN "00000000000000000000000000000101" => fio_result <= "00000010000000000000010100010011";
					WHEN "00000000000000000000000000000110" => fio_result <= "00000010000100000000010100010011";
					WHEN "00000000000000000000000000000111" => fio_result <= "00000010001000000000010100010011";
					WHEN "00000000000000000000000000001000" => fio_result <= "00000010001100000000010100010011";
					WHEN "00000000000000000000000000001001" => fio_result <= "00000010010000000000010100010011";
					WHEN "00000000000000000000000000001010" => fio_result <= "00000000011100000000011100010011";
					WHEN "00000000000000000000000000001011" => fio_result <= "11111101010111111111000011101111";
					WHEN "00000000000000000000000000001100" => fio_result <= "00000001010000000000010100010011";
					WHEN "00000000000000000000000000001101" => fio_result <= "00000000011100000000011010010011";
					WHEN "00000000000000000000000000001110" => fio_result <= "00000010110101110000010001100011";
					WHEN "00000000000000000000000000001111" => fio_result <= "00000000000000000000000000000000";
					when others => report "unreachable" severity failure;
				END CASE;
		END PROCESS;
		
END ARCHITECTURE;