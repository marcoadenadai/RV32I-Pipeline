LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE ADDER_PACKAGE IS
   COMPONENT ADDER
   PORT (
		A	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		S 	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
   );
   END COMPONENT;
END ADDER_PACKAGE; 