LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE BRANCH_COMPARE_PACKAGE IS
   COMPONENT BRANCH_COMPARE 
   PORT (
      clock    				: IN STD_LOGIC := '0';
		Reset						: IN STD_LOGIC := '0';
		BRANCH_OP				: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		REG_1_IN       		: IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
		REG_2_IN       		: IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
      DECISION       : OUT STD_LOGIC
	);
   END COMPONENT;
END BRANCH_COMPARE_PACKAGE;