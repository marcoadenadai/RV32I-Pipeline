LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;

ENTITY AND_BRANCH IS
   PORT (
		BRANCH_DO_IT            : IN STD_LOGIC;
		COMPARE_BRANCH_OUT		: IN STD_LOGIC;
		AND_OUT	: OUT STD_LOGIC
		);
END ENTITY;

ARCHITECTURE AND_BRANCH_Arch OF AND_BRANCH IS
	
	BEGIN

        AND_OUT <= BRANCH_DO_IT AND COMPARE_BRANCH_OUT; 
		
END ARCHITECTURE;