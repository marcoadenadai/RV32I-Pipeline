
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;
USE ieee.std_logic_signed.all;

LIBRARY work;
USE work.PC_PACKAGE.all;

USE work.ROM_PACKAGE.all;

USE work.REGPIPE_IF_DF_PACKAGE.all;

USE work.BancoRegistradores_PACKAGE.all;

USE work.REGPIPE_ID_EX_PACKAGE.all;

USE work.BRANCH_COMPARE_PACKAGE.all;

USE work.MUX_ALU_1_PACKAGE.all;

USE work.MUX_ALU_2_PACKAGE.all;

USE work.ULA_PACKAGE.all;

USE work.IMM_HANDLER_PACKAGE.all;

USE work.REGPIPE_EX_MEM_PACKAGE.all;

USE work.AND_BRANCH_PACKAGE.all;

USE work.RAM_PACKAGE.all;

USE work.REGPIPE_MEM_WB_PACKAGE.all;

USE work.MUX_MEM_TO_REG_PACKAGE.all;


ENTITY PROCESSADOR IS
	PORT(
		CLK : IN STD_LOGIC;
		RESET: IN STD_LOGIC;
		
		--CONTROLE-----------------------
		REGWRITE: IN STD_LOGIC;
		BRANCH_OP: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		MEM_WRITE: IN STD_LOGIC;
		MEM_READ: IN STD_LOGIC
		
		--Saida_PC : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		--Saida_ROM : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		--Saida_TEST : OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
	);

END ENTITY;

ARCHITECTURE PROCESSADOR_ARCH OF PROCESSADOR IS
	--variable PC_IN: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL PC_OUT: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL PC_NEXT: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ROM_INSTRUCTION: STD_LOGIC_VECTOR(31 DOWNTO 0);


--	SIGNAL ROM_INSTRUCTION: STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
--	--SIGNAL TEST_RETURN: STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
	SIGNAL REGPIPE_IF_DF_SAIDA_PC:  STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000"; --Serão as entrada do estágio de DF
	SIGNAL REGPIPE_IF_DF_SAIDA_INSTRUCTION:  STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";--Serão as entrada do estágio de DF
--	
	SIGNAL myCLK: STD_LOGIC;
	SIGNAL myRESET: STD_LOGIC;
	SIGNAL myREGWRITE: STD_LOGIC;
	SIGNAL myBRANCH_OP: STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL myMEM_READ: STD_LOGIC;
	SIGNAL myMEM_WRITE: STD_LOGIC;
	
	SIGNAL REG_OUT_1: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL REG_OUT_2: STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	SIGNAL REGPIPE_ID_EX_SAIDA_PC: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL REGPIPE_ID_EX_SAIDA_REG_OUT_1: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL REGPIPE_ID_EX_SAIDA_REG_OUT_2: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL REGPIPE_ID_EX_SAIDA_INSTRUCTION:  STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	SIGNAL DECISION_BRANCH_OUT: STD_LOGIC;
	SIGNAL MUX_OUT_EM_1:  STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL MUX_OUT_EM_2:  STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	SIGNAL ULA_RESULT:  STD_LOGIC_VECTOR(31 DOWNTO 0);
	
	SIGNAL IMM_HANDLER_OUT: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL RD_HANDLER_OUT: STD_LOGIC_VECTOR(4 DOWNTO 0);
	
	SIGNAL REGPIPE_EX_MEM_SAIDA_PC: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL REGPIPE_EX_MEM_SAIDA_BRANCH_CONTROL: STD_LOGIC;
	SIGNAL REGPIPE_EX_MEM_SAIDA_ULA: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL REGPIPE_EX_MEM_SAIDA_REG_OUT_2: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL REGPIPE_EX_MEM_SAIDA_RD_HANDLER_2: STD_LOGIC_VECTOR(4 DOWNTO 0);
	
	SIGNAL AND_BRANCH_OUT: STD_LOGIC;
	SIGNAL RAM_OUT: STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL AUX_UNSIGNED: UNSIGNED(31 DOWNTO 0);
	
	SIGNAL REGPIPE_MEM_WB_SAIDA_PC, REGPIPE_MEM_WB_SAIDA_RAM_OUT, REGPIPE_MEM_WB_SAIDA_ULA :STD_LOGIC_VECTOR(31 DOWNTO 0); 
	SIGNAL REGPIPE_MEM_WB_SAIDA_RD_HANDLER : STD_LOGIC_VECTOR(4 DOWNTO 0); 
	
	SIGNAL MUX_MEM_TO_REG_SAIDA: STD_LOGIC_VECTOR(31 DOWNTO 0);
	
 BEGIN
	
	myCLK <= CLK;
	myRESET <= RESET;
	myREGWRITE <= REGWRITE;
	myBRANCH_OP <= BRANCH_OP;
	myMEM_WRITE <= MEM_WRITE;
	myMEM_READ <= MEM_READ;
   ------------------------------------ IF ---------------------------------------
	--ADICONAR PC_MUX (PRONTO)
	
	PC_C0: PC PORT MAP(myCLK, myRESET, PC_NEXT, PC_OUT, PC_NEXT);
	ROM_C1: ROM PORT MAP(myCLK, myRESET, PC_OUT, ROM_INSTRUCTION);
	
	REGPIPE_IF_DF_C3: REGPIPE_IF_DF PORT MAP(myCLK, myRESET, PC_OUT, REGPIPE_IF_DF_SAIDA_PC, ROM_INSTRUCTION, REGPIPE_IF_DF_SAIDA_INSTRUCTION);
	
	------------------------------------ DF ---------------------------------------
	
	BANCO_REG: BancoRegistradores PORT MAP(myREGWRITE, myCLK, myRESET, "00000", "00001", "00001", "11111111111111111111111111111111",REG_OUT_1, REG_OUT_2);
	
	REGPIPE_ID_EX_C4: REGPIPE_ID_EX PORT MAP(myCLK, myRESET, REGPIPE_IF_DF_SAIDA_PC, REGPIPE_ID_EX_SAIDA_PC , REG_OUT_1, REGPIPE_ID_EX_SAIDA_REG_OUT_1, REG_OUT_2, REGPIPE_ID_EX_SAIDA_REG_OUT_2, REGPIPE_IF_DF_SAIDA_INSTRUCTION, REGPIPE_ID_EX_SAIDA_INSTRUCTION);
	
	------------------------------------ EX ----------------------------------------
	
	BRANCH_COMPARE_c5: BRANCH_COMPARE PORT MAP(myCLK, myRESET, myBRANCH_OP, REGPIPE_ID_EX_SAIDA_REG_OUT_1, REGPIPE_ID_EX_SAIDA_REG_OUT_2, DECISION_BRANCH_OUT);
	--ESTA SAINDO SINAL ERRADO (VER)
	
	
	
	MUX_ALU_1_C6: MUX_ALU_1 PORT MAP('0', REGPIPE_ID_EX_SAIDA_PC, REGPIPE_ID_EX_SAIDA_REG_OUT_1, MUX_OUT_EM_1); -- BRANCH_DO_IT, PC_IN_MUX, REG_OUT_1, MUX_OUT_ALU_1(SAIDA)
	
	MUX_ALU_2_C7: MUX_ALU_2 PORT MAP('0', "00000000000000000000000000000000", REGPIPE_ID_EX_SAIDA_REG_OUT_2, MUX_OUT_EM_2);-- ALU_SRC, IMM, REG_OUT_2, MUX_OUT_ALU_2(SAIDA)
	
	ULA_C8: ULA PORT MAP(myCLK, myRESET, "0010", MUX_OUT_EM_1, MUX_OUT_EM_2, ULA_RESULT); --CLOCK, RESET, ALUOP, A, B, ULAOUT
	
	--ADICIONAR IMM. HANDLER (PRONTO) (N TA FUNCIONANDO)
	IMM_HANDLER_C9: IMM_HANDLER PORT MAP("011", REGPIPE_ID_EX_SAIDA_INSTRUCTION, RD_HANDLER_OUT, IMM_HANDLER_OUT); -- IMM_TYPE, INSTRUCTION, RD(SAIDA), IMM_OUT(SAIDA)	
	
	
	--ADICIONAR REGPIPE_EX_MEM (PRONTO)
	REGPIPE_EX_MEM_C10: REGPIPE_EX_MEM PORT MAP(myCLK, myRESET, REGPIPE_ID_EX_SAIDA_PC, REGPIPE_EX_MEM_SAIDA_PC, DECISION_BRANCH_OUT, REGPIPE_EX_MEM_SAIDA_BRANCH_CONTROL,ULA_RESULT, REGPIPE_EX_MEM_SAIDA_ULA, REGPIPE_ID_EX_SAIDA_REG_OUT_2, REGPIPE_EX_MEM_SAIDA_REG_OUT_2, RD_HANDLER_OUT, REGPIPE_EX_MEM_SAIDA_RD_HANDLER_2);--CLOCK, RESET, PCIN, PCOUT, BRANCH_COMPARE_IN, BRANCH_COMPARE_OUT, ALU_IN, ALU_OUT, REG_IN, REG_OUT, RD_IN, RD_OUT
	
	------------------------------------- MEM -------------------------------------

	
	--ADICIONAR PORTA AND (PRONTO)
	AND_BRANCH_C11: AND_BRANCH PORT MAP('1', REGPIPE_EX_MEM_SAIDA_BRANCH_CONTROL, AND_BRANCH_OUT); --BRANCH_DO_IT, COMPARE_BRANCH_OUT, AND_OUT(SAIDA)
	
	
	--ADICIONAR RAM (PRONTO)
	AUX_UNSIGNED <= UNSIGNED(REGPIPE_EX_MEM_SAIDA_ULA);

	RAM_C12: RAM PORT MAP(myCLK, myRESET, myMEM_WRITE, myMEM_READ, AUX_UNSIGNED, REGPIPE_EX_MEM_SAIDA_REG_OUT_2, RAM_OUT);--CLOCK,RESET, MEM_WRITE, MEM_READ, ADDR, WRITE_DATA, MEM_OUT
	
	--ADICIONAR REGPIPE_MEM_WB (PRONTO)
	REGPIPE_MEM_WB_C13: REGPIPE_MEM_WB PORT MAP(myCLK, myRESET, REGPIPE_EX_MEM_SAIDA_PC, REGPIPE_MEM_WB_SAIDA_PC, RAM_OUT, REGPIPE_MEM_WB_SAIDA_RAM_OUT, REGPIPE_EX_MEM_SAIDA_ULA, REGPIPE_MEM_WB_SAIDA_ULA, REGPIPE_EX_MEM_SAIDA_RD_HANDLER_2, REGPIPE_MEM_WB_SAIDA_RD_HANDLER); --clock, reset, PCIN, PC_OUT, MEM_IN, MEM_OUT, ALU_IN, ALU_OUT, RD_IN, RD_OUT

	
	------------------------------------- WB ---------------------------------------
	--ADICIONAR MUX WB 3X1 (PRONTO)
	MUX_MEM_TO_REG_C14: MUX_MEM_TO_REG PORT MAP("00", REGPIPE_MEM_WB_SAIDA_RAM_OUT, REGPIPE_MEM_WB_SAIDA_ULA, REGPIPE_MEM_WB_SAIDA_PC, MUX_MEM_TO_REG_SAIDA);--MEM_TO_REG, OUT_MEMORY, ALU_RESULT, PC_OUT, MUX_OUT_MEM_TO_REG(SAIDA)
	
	
--FALTA OS REGISTRADORES DE PIPE DOS SINAIS(ADICIONAR DENTRO DOS OUTROS REG DE PIPE)

--TEM UM ERRO NA SIMULA'C~AO, OBSERVAR LA QUAL O ERRO E CORRIGIR 





	--------------------------------------------------------------------------------

	
--	ROM_C1: ROM PORT MAP(PC_VALUE, ROM_INSTRUCTION, myCLK, myRESET);
--	
   
--	
--	Saida_TEST <= REGPIPE_IF_DF_SAIDA_INSTRUCTION;
--	Saida_PC <= PC_VALUE;
--	Saida_ROM <= ROM_INSTRUCTION;
	
END ARCHITECTURE;