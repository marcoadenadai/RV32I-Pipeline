LIBRARY ieee;
USE ieee.std_logic_1164.all;
LIBRARY work;
USE work.ROM_PACKAGE.all;
USE work.PC_PACKAGE.all;
USE work.ADDER_PACKAGE.all;

ENTITY PROCESSADOR_tb IS
END ENTITY;


ARCHITECTURE PROCESSADOR_tb_arch OF PROCESSADOR_tb IS
	constant PERIODO : time := 10 ns;

	SIGNAL CLK : STD_LOGIC := '0';
	SIGNAL RESET: STD_LOGIC;
	SIGNAL PC : STD_LOGIC_VECTOR(31 DOWNTO 0);
	SIGNAL ROM : STD_LOGIC_VECTOR(31 DOWNTO 0);
BEGIN
	--C0_PC : PC PORT MAP(myCLK, myRESET, PC2_VALUE, PC_VALUE);
	CLK <= NOT CLK after PERIODO/2;
 
 
END ARCHITECTURE;