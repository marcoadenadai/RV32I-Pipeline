LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE REGPIPE_MEM_WB_PACKAGE IS
   COMPONENT REGPIPE_MEM_WB
      PORT (
			clock    				: IN STD_LOGIC := '0';
			Reset						: IN STD_LOGIC := '0';
			
			PCIn						: IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
			PCOut        			: OUT STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
			
			MEM_IN					: IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
			MEM_OUT       			: OUT STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
			
			ALU_IN					: IN STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
			ALU_OUT       			: OUT STD_LOGIC_VECTOR(31 DOWNTO 0) := "00000000000000000000000000000000";
			
			RD_IN						: IN STD_LOGIC_VECTOR(4 DOWNTO 0) := "00000";
			RD_OUT       			: OUT STD_LOGIC_VECTOR(4 DOWNTO 0) := "00000";
			
			ctl_RegWrite_IN		: IN STD_LOGIC := '0';
			ctl_RegWrite_OUT		: OUT STD_LOGIC := '0';
			
			ctl_MemToReg_IN		: IN STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
			ctl_MemToReg_OUT		: OUT STD_LOGIC_VECTOR(1 DOWNTO 0) := "00"
		);
   END COMPONENT;
END REGPIPE_MEM_WB_PACKAGE;