LIBRARY ieee;
USE ieee.std_logic_1164.all;

PACKAGE ULA_PACKAGE IS
   COMPONENT ULA
      PORT(
			ULAop			:IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
			A, B			:IN	STD_LOGIC_VECTOR(31 DOWNTO 0);
			ULAout 			:OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
		);
   END COMPONENT;
END ULA_PACKAGE;